//--------------------------------------
//-- debugCode.v
//--
//-- This file provides a way to add code to
//-- the simulation. Examples are given below.
//-- Uncomment the parts you want to have included
//-- in a.out when you compile your top-level cell,
//--
//--     0_LC4_Top{sch}
//--
//-- (Note: There is an  `include "debugCode.v"
//-- compiler directive in that cell's verilog code.)
//------------------------------------

// always @(PCout) begin
//     #1 $display("(t=%0d)    PCout=%b  "         , ($time-1),  PCout);
// end
// always @(PCout) begin
//     #1 $display("(t=%0d)    PCout=%h  "         , ($time-1),  PCout);
// end
// always @(PCmux) begin
//     #1 $display("(t=%0d)    PCmux=%b  "         , ($time-1),  PCmux);
// end
// always @(nextPC) begin
//     #1 $display("(t=%0d)    nextPC=%h  "         , ($time-1),  nextPC);
// end
 always @(IR) begin
     #1 $display("(t=%0d)    IR[15:12]=%b "      , ($time-1),  IR[15:12] );
        $display("(t=%0d)    IR[11:8] =%b "      , ($time-1),  IR[11:9]  );
        $display("(t=%0d)    IR[8:6]  =%b "      , ($time-1),  IR[8:6]   );
        $display("(t=%0d)    IR[5:3]  =%b "      , ($time-1),  IR[5:3]   );
        $display("(t=%0d)    IR[2:0]  =%b "      , ($time-1),  IR[2:0]   );
 end
// always @(IR[8:0]) begin
//     #1 $display("(t=%0d)    IR[8:0]=%b "        , ($time-1),  IR[8:0]);
// end
 always @ ( Rwe ) begin
     #1 $display("(t=%0d)    Rwe=%b "            , ($time-1),  Rwe);
 end
 always @ ( PipeRwe ) begin
     #1 $display("(t=%0d)    PipeRwe=%b "            , ($time-1),  PipeRwe);
 end
 always @ ( DRmux ) begin
     #1 $display("(t=%0d)    DRmux=%b "          , ($time-1),  DRmux);
 end
 always @ ( DR ) begin
     #1 $display("(t=%0d)    DR=%b "             , ($time-1),  DR[2:0]);
 end
// always @ ( out1 ) begin
//     #1 $display("(t=%0d)    out1=%b "           , ($time-1),  out1);
// end
// always @ ( out2 ) begin
//     #1 $display("(t=%0d)    out2=%b "           , ($time-1),  out2);
// end
// always @ ( ALUout ) begin
//     #1 $display("(t=%0d)    ALUout=%b "         , ($time-1),  ALU.out);
// end
// always @ ( immed ) begin
//     #1 $display("(t=%0d)    immed=%b "          , ($time-1),  immed);
// end
// always @ ( DMEMout ) begin
//     #1 $display("(t=%0d)    DMEMout=%b "        , ($time-1),  DMEMout);
// end
// always @ ( PipeINmux ) begin
//     #1 $display("(t=%0d)    PipeINmux=%b "          , ($time-1),  PipeINmux);
// end

 always @ ( Mwe ) begin
     #1 $display("(t=%0d)    Mwe=%b "            , ($time-1),  Mwe);
 end
 always @ ( PipeMwe ) begin
     #1 $display("(t=%0d)    PipeMwe=%b "            , ($time-1),  PipeMwe);
 end
// always @ ( BR ) begin
//     #1 $display("(t=%0d)    BR=%b "             , ($time-1),  BR);
// end
// always @ ( I_interface ) begin
//     #1 $display("(t=%0d)    I_interface=[ %b ] ", ($time-1),  I_interface);
// end
// always @ ( D_interface ) begin
//     #1 $display("(t=%0d)    D_interface=[ %b ] ", ($time-1),  D_interface);
// end
 always @ ( ALUsel1 ) begin
     #1 $display("(t=%0d)    ALUsel1=%b "            , ($time-1),  ALUsel1);
 end

 always @ ( ALUsel2 ) begin
     #1 $display("(t=%0d)    ALUsel2=%b "            , ($time-1),  ALUsel2);
 end

 always @ ( ALUinput1 ) begin
     #1 $display("(t=%0d)    ALUInput1=%b "            , ($time-1),  ALUinput1);
 end

 always @ ( ALUinput2 ) begin
     #1 $display("(t=%0d)    ALUInput2=%b "            , ($time-1),  ALUinput2);
 end
 always @ ( reg_in ) begin
     #1 $display("(t=%0d)    reg_in=%b "         , ($time-1),  reg_in);
 end
 always @ ( out1 ) begin
     #1 $display("(t=%0d)    out1=%b "         , ($time-1),  out1);
 end
 always @ ( out2 ) begin
     #1 $display("(t=%0d)    out2=%b "         , ($time-1),  out2);
 end
 always @ ( ALUsel1 ) begin
    #1 $display("(t=%0d)    ALUsel1=%b "         , ($time-1),  ALUsel1);
 end
 always @ ( ALUsel2 ) begin
    #1 $display("(t=%0d)    ALUsel2=%b "         , ($time-1),  ALUsel2);
 end
